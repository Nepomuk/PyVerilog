
module TOP( in, out );
input  in;
output  out;
INVD1 U0( .I( in ), .ZN( out ) );
endmodule
